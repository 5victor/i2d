/* generator.sv
 *
 * Copyright Victor Wen, vic7tor@gmail.com
 * This code publish under GNU GPL License
 *
 * Description:
 *
 * TODO
 */

`include "i2d_core_defines.sv"

class generator;
rand instr_t instr;

function void post_randomize();

endfunction
endclass
